interface interfejs (
 input bit clk
);

logic rst_n;
logic in;
logic out;

endinterface
